module Grey_Square (
    output P,H,
    input A,B
);

or Prop (P,A,B);
xor Gen (H,A,B);

endmodule